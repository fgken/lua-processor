module cpu(clk);
	input wire clk;

	// Fetch
	
	// Decode
	
	// Execute
	
	// Memory access

	// Write Back

endmodule
